
-- Buffer Testbench -- 									

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;


entity buffertb is 

end entity;



architecture buffertbarc is 

begin 


end buffertbarc;










-- Buffer Testbench Plan --

-- Generate input 
-- Gneerate clock 
	-- Make it run at 1Khz.
-- Send said input to the array 
	-- 1024 values 
	-- Once full send those bits to the output CALC
-- Empty array to an output
-- 